netcdf new {
dimensions:
	x    = 2;
	y    = 3;
	time = UNLIMITED ; // (12 currently)
variables:
        float a(x,y);
	int date(time) ;
	int time(time) ;
        short b(time, y, x);
data:
 a = 1.0, 2.0, 3.0, 4.0, 5.0, 6.0;

 date = 840116, 840214, 840316, 840415, 840516, 840615, 840716, 840816, 
    840915, 841016, 841115, 841216 ;

 time = 1, 2, 3, 4, 5, 6, 7, 8, 9, 10, 11, 12 ;
  
 b = 1, 1, 2, 2, 3, 3,
     4, 4, 5, 5, 6, 6,
     7, 7, 8, 8, 9, 9,
    10, 10, 11, 11, 12, 12,
    13, 13, 14, 14, 15, 15,
    16, 16, 17, 17, 18, 18,
    19, 19, 20, 20, 21, 22,
    23, 23, 24, 24, 25, 25,
    26, 26, 27, 27, 28, 28,
    29, 29, 30, 30, 31, 31,
    32, 32, 33, 33, 34, 34,
    35, 35, 36, 36, 37, 37 ;
}
